module ENCODER83_TB();

reg  [7:0] X;
wire [2:0] Y;

encoder83 DUT(.x(X), .y(Y));

initial
begin
    #10 X=8'b00000000;
    #10 X=8'b00000001;
    #10 X=8'b00000010;
    #10 X=8'b00000100;
    #10 X=8'b00001000;
    #10 X=8'b00010000;
    #10 X=8'b00100000;
    #10 X=8'b01000000;
    #10 X=8'b10000000;
    #10 X=8'b01000100;
    #10 X=8'b00000011;
    #10 X=8'b00000001;
    #10
    $finish;
end

endmodule
